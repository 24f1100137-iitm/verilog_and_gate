# And_gate design.sv in EDA playground
// Code your design here
module And(
  input wire x,y,
  output wire z
);
  assign z=x&y; // assign the value of x and y in z //
endmodule
